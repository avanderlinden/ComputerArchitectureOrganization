library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memory is
	port
	(
		clk			: in  std_logic;
		rst			: in  std_logic;
		memread			: in  std_logic;
		memwrite		: in  std_logic;
		address1		: in  std_logic_vector (31 downto 0);
		address2		: in  std_logic_vector (31 downto 0);
		writedata		: in  std_logic_vector (31 downto 0);
		instruction		: out std_logic_vector (31 downto 0);
		readdata		: out std_logic_vector (31 downto 0)
	);
end memory;

architecture behavior of memory is
	type ramcell is array (0 to 255) of std_logic_vector (7 downto 0);
	signal ram			: ramcell;
	signal masked1, masked2		: std_logic_vector (7 downto 0);
	signal selector1, selector2	: natural range 0 to 255;
begin
	masked1 <= address1 (7 downto 2) & "00";
	masked2 <= address2 (7 downto 2) & "00";
	selector1 <= to_integer (unsigned (masked1));
	selector2 <= to_integer (unsigned (masked2));

	process (clk, rst, memread, memwrite, address1, address2, writedata)
	begin
		if (rising_edge (clk)) then
			if (rst = '1') then
				ram (  0) <= "11111111"; -- lui	$0,-1
				ram (  1) <= "11111111";
				ram (  2) <= "00000000";
				ram (  3) <= "00111100";
				ram (  4) <= "11111111"; -- lui	$1,-1
				ram (  5) <= "11111111";
				ram (  6) <= "00000001";
				ram (  7) <= "00111100";
				ram (  8) <= "11111111"; -- ori	$1,$1,-1
				ram (  9) <= "11111111";
				ram ( 10) <= "00100001";
				ram ( 11) <= "00110100";
				ram ( 12) <= "00110000"; -- addi	$1,$0,48
				ram ( 13) <= "00000000";
				ram ( 14) <= "00000001";
				ram ( 15) <= "00100000";
				ram ( 16) <= "01000010"; -- srl 	$1,$1,1
				ram ( 17) <= "00001000";
				ram ( 18) <= "00000001";
				ram ( 19) <= "00000000";
				ram ( 20) <= "01000011"; -- sra 	$1,$1,1
				ram ( 21) <= "00001000";
				ram ( 22) <= "00000001";
				ram ( 23) <= "00000000";
				ram ( 24) <= "11101000"; -- addiu	$1,$1,-24
				ram ( 25) <= "11111111";
				ram ( 26) <= "00100001";
				ram ( 27) <= "00100100";
				ram ( 28) <= "01000011"; -- sra	$1,$1,1
				ram ( 29) <= "00001000";
				ram ( 30) <= "00000001";
				ram ( 31) <= "00000000";
				ram ( 32) <= "00001010"; -- j	B
				ram ( 33) <= "00000000";
				ram ( 34) <= "00000000";
				ram ( 35) <= "00001000";
				ram ( 36) <= "00000001"; -- lui	$2,1
				ram ( 37) <= "00000000";
				ram ( 38) <= "00000010";
				ram ( 39) <= "00111100";
				ram ( 40) <= "00101010"; -- addi	$3,$0,42
				ram ( 41) <= "00000000";
				ram ( 42) <= "00000011";
				ram ( 43) <= "00100000";
				ram ( 44) <= "11111010"; -- addiu	$4,$3,-6
				ram ( 45) <= "11111111";
				ram ( 46) <= "01100100";
				ram ( 47) <= "00100100";
				ram ( 48) <= "00001010"; -- jal	B
				ram ( 49) <= "00000000";
				ram ( 50) <= "00000000";
				ram ( 51) <= "00001100";
				ram ( 52) <= "00001101"; -- j	C
				ram ( 53) <= "00000000";
				ram ( 54) <= "00000000";
				ram ( 55) <= "00001000";
				ram ( 56) <= "00100000"; -- add	$5,$4,$3
				ram ( 57) <= "00101000";
				ram ( 58) <= "10000011";
				ram ( 59) <= "00000000";
				ram ( 60) <= "00100001"; -- addu	$6,$5,$5
				ram ( 61) <= "00110000";
				ram ( 62) <= "10100101";
				ram ( 63) <= "00000000";
				ram ( 64) <= "00100100"; -- and	$7,$6,$3
				ram ( 65) <= "00111000";
				ram ( 66) <= "11000011";
				ram ( 67) <= "00000000";
				ram ( 68) <= "11101001"; -- andi	$8,$1,-23
				ram ( 69) <= "11111111";
				ram ( 70) <= "00101000";
				ram ( 71) <= "00110000";
				ram ( 72) <= "00100111"; -- nor	$9,$8,$6
				ram ( 73) <= "01001000";
				ram ( 74) <= "00000110";
				ram ( 75) <= "00000001";
				ram ( 76) <= "00100101"; -- or	$10,$9,$5
				ram ( 77) <= "01010000";
				ram ( 78) <= "00100101";
				ram ( 79) <= "00000001";
				ram ( 80) <= "00000010"; -- srl	$11,$10,8
				ram ( 81) <= "01011010";
				ram ( 82) <= "00001010";
				ram ( 83) <= "00000000";
				ram ( 84) <= "00000000"; -- sll	$12,$11,4
				ram ( 85) <= "01100001";
				ram ( 86) <= "00001011";
				ram ( 87) <= "00000000";
				ram ( 88) <= "00100010"; -- sub	$13,$12,$3
				ram ( 89) <= "01101000";
				ram ( 90) <= "10000011";
				ram ( 91) <= "00000001";
				ram ( 92) <= "00100011"; -- subu	$14,$12,$13
				ram ( 93) <= "01110000";
				ram ( 94) <= "10001101";
				ram ( 95) <= "00000001";
				ram ( 96) <= "00000111"; -- xori	$15,$14,7
				ram ( 97) <= "00000000";
				ram ( 98) <= "11001111";
				ram ( 99) <= "00111001";
				ram (100) <= "00100110"; -- xor	$16,$15,$14
				ram (101) <= "10000000";
				ram (102) <= "11101110";
				ram (103) <= "00000001";
				ram (104) <= "11111111"; -- beq	$14,$5,D
				ram (105) <= "11111111";
				ram (106) <= "11000101";
				ram (107) <= "00010001";
				ram (108) <= "00000001"; -- beq	$14,$3,F
				ram (109) <= "00000000";
				ram (110) <= "11000011";
				ram (111) <= "00010001";
				ram (112) <= "00011100"; -- j	E
				ram (113) <= "00000000";
				ram (114) <= "00000000";
				ram (115) <= "00001000";
				ram (116) <= "00000001"; -- bne	$4,$5,H
				ram (117) <= "00000000";
				ram (118) <= "10000101";
				ram (119) <= "00010100";
				ram (120) <= "00011110"; -- j	G
				ram (121) <= "00000000";
				ram (122) <= "00000000";
				ram (123) <= "00001000";
				ram (124) <= "11111111"; -- bne	$3,$14,H
				ram (125) <= "11111111";
				ram (126) <= "01101110";
				ram (127) <= "00010100";
				ram (128) <= "00000001"; -- bgez	$0,J
				ram (129) <= "00000000";
				ram (130) <= "00000001";
				ram (131) <= "00000100";
				ram (132) <= "00100001"; -- j	I
				ram (133) <= "00000000";
				ram (134) <= "00000000";
				ram (135) <= "00001000";
				ram (136) <= "11111111"; -- bgez	$1,J
				ram (137) <= "11111111";
				ram (138) <= "00100001";
				ram (139) <= "00000100";
				ram (140) <= "00000001"; -- bgez	$3,L
				ram (141) <= "00000000";
				ram (142) <= "01100001";
				ram (143) <= "00000100";
				ram (144) <= "00100100"; -- j	K
				ram (145) <= "00000000";
				ram (146) <= "00000000";
				ram (147) <= "00001000";
				ram (148) <= "11111111"; -- bgtz	$0,L
				ram (149) <= "11111111";
				ram (150) <= "00000000";
				ram (151) <= "00011100";
				ram (152) <= "11111111"; -- bgtz	$1,M
				ram (153) <= "11111111";
				ram (154) <= "00100000";
				ram (155) <= "00011100";
				ram (156) <= "00000001"; -- bgtz	$3,O
				ram (157) <= "00000000";
				ram (158) <= "01100000";
				ram (159) <= "00011100";
				ram (160) <= "00101000"; -- j	N
				ram (161) <= "00000000";
				ram (162) <= "00000000";
				ram (163) <= "00001000";
				ram (164) <= "00000001"; -- blez	$0,Q
				ram (165) <= "00000000";
				ram (166) <= "00000000";
				ram (167) <= "00011000";
				ram (168) <= "00101010"; -- j	P
				ram (169) <= "00000000";
				ram (170) <= "00000000";
				ram (171) <= "00001000";
				ram (172) <= "11111111"; -- blez	$3,Q
				ram (173) <= "11111111";
				ram (174) <= "01100000";
				ram (175) <= "00011000";
				ram (176) <= "00000001"; -- blez	$1,S
				ram (177) <= "00000000";
				ram (178) <= "00100000";
				ram (179) <= "00011000";
				ram (180) <= "00101101"; -- j	R
				ram (181) <= "00000000";
				ram (182) <= "00000000";
				ram (183) <= "00001000";
				ram (184) <= "11111111"; -- bltz	$0,S
				ram (185) <= "11111111";
				ram (186) <= "00000000";
				ram (187) <= "00000100";
				ram (188) <= "11111111"; -- bltz	$3,T
				ram (189) <= "11111111";
				ram (190) <= "01100000";
				ram (191) <= "00000100";
				ram (192) <= "00000001"; -- bltz	$1,V
				ram (193) <= "00000000";
				ram (194) <= "00100000";
				ram (195) <= "00000100";
				ram (196) <= "00110001"; -- j	U
				ram (197) <= "00000000";
				ram (198) <= "00000000";
				ram (199) <= "00001000";
				ram (200) <= "11111000"; -- addi	$17,$0,248
				ram (201) <= "00000000";
				ram (202) <= "00010001";
				ram (203) <= "00100000";
				ram (204) <= "11111100"; -- sw	$1,-4($17)
				ram (205) <= "11111111";
				ram (206) <= "00100001";
				ram (207) <= "10101110";
				ram (208) <= "00000000"; -- sw	$3,0($17)
				ram (209) <= "00000000";
				ram (210) <= "00100011";
				ram (211) <= "10101110";
				ram (212) <= "00000100"; -- sw	$4,4($17)
				ram (213) <= "00000000";
				ram (214) <= "00100100";
				ram (215) <= "10101110";
				ram (216) <= "00111001"; -- j	X
				ram (217) <= "00000000";
				ram (218) <= "00000000";
				ram (219) <= "00001000";
				ram (220) <= "11111000"; -- addi	$17,$17,-8
				ram (221) <= "11111111";
				ram (222) <= "00110001";
				ram (223) <= "00100010";
				ram (224) <= "00111100"; -- j	Y
				ram (225) <= "00000000";
				ram (226) <= "00000000";
				ram (227) <= "00001000";
				ram (228) <= "11111100"; -- lw	$18,-4($17)
				ram (229) <= "11111111";
				ram (230) <= "00110010";
				ram (231) <= "10001110";
				ram (232) <= "00000000"; -- lw	$19,0($17)
				ram (233) <= "00000000";
				ram (234) <= "00110011";
				ram (235) <= "10001110";
				ram (236) <= "00110111"; -- j	W
				ram (237) <= "00000000";
				ram (238) <= "00000000";
				ram (239) <= "00001000";
				ram (240) <= "00001100"; -- lw	$20,12($17)
				ram (241) <= "00000000";
				ram (242) <= "00110100";
				ram (243) <= "10001110";
				ram (244) <= "00111101"; -- j	Z
				ram (245) <= "00000000";
				ram (246) <= "00000000";
				ram (247) <= "00001000";
				for i in 248 to 255 loop
					ram (i) <= std_logic_vector (to_unsigned (0, 8));
				end loop;
			else
				if (memwrite = '1') then
					ram (selector2 + 0) <= writedata (7 downto 0);
					ram (selector2 + 1) <= writedata (15 downto 8);
					ram (selector2 + 2) <= writedata (23 downto 16);
					ram (selector2 + 3) <= writedata (31 downto 24);
				end if;
			end if;
		end if;
	end process;
	instruction <= ram (selector1 + 3) & ram (selector1 + 2) & ram (selector1 + 1) & ram (selector1 + 0);
	with memread select
		readdata <=	std_logic_vector (to_unsigned (0, 32)) when '0',
				ram (selector2 + 3) & ram (selector2 + 2) & ram (selector2 + 1) & ram (selector2 + 0) when others;
end behavior;
